module hello (A, B); //Module named hello, define inputs and outputs

    input A; //declare input
    output B;//declare output


    assign B = A;

endmodule